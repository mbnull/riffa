`ifndef GOWIN_VH
`define GOWIN_VH 1



`endif
